// femtorv32, a minimalistic RISC-V RV32I core
//    (minus SYSTEM and FENCE that are not implemented)
//
//       Bruno Levy, May-June 2020
//
// This file: the "System on Chip" that goes with femtorv32.

/*************************************************************************************/


`default_nettype none // Makes it easier to detect typos !


/*************************************************************************************/

`define NRV_FREQ 50 // Base frequency in MHz

`ifndef NRV_RESET_ADDR
   `define NRV_RESET_ADDR 0
`endif

`ifndef NRV_ADDR_WIDTH
   `define NRV_ADDR_WIDTH 24
`endif

`ifndef NRV_RAM_SIZE
   `define NRV_RAM_SIZE 64 * 1024
`endif

`define NRV_IO_BUTTONS
`define NRV_IO_LEDS
`define NRV_IO_UART
`define NRV_IO_HARDWARE_CONFIG

/*************************************************************************************/

module femtosoc (
   input  wire       pclk
  ,input  wire       RESET
  ,output wire       D1, D2, D3, D4, D5
  ,input  wire       RXD
  ,output wire       TXD
  ,input  wire [5:0] buttons
);


  wire clk;

  femtoPLL #(
     .freq(`NRV_FREQ)
  ) pll (
      .pclk(pclk)
     ,.clk(clk)
  );

   reg [15:0] reset_cnt = 0;
   wire       reset = &(reset_cnt);

/* verilator lint_off WIDTH */   
`ifdef NRV_NEGATIVE_RESET
   always @(posedge clk,negedge RESET) begin
      if(!RESET) begin
         reset_cnt <= 0;
      end else begin
         reset_cnt <= reset_cnt + !reset;
      end
   end
`else
   always @(posedge clk,posedge RESET) begin
      if(RESET) begin
         reset_cnt <= 0;
      end else begin
         reset_cnt <= reset_cnt + !reset;
      end
   end
`endif
/* verilator lint_on WIDTH */   
   
/***************************************************************************************************
 *
 * Memory and memory interface
 * memory map:
 *   address[21:2] RAM word address (4 Mb max).
 *   address[23:22]   00: RAM
 *                    01: IO page (1-hot)  (starts at 0x400000)
 *                    10: SPI Flash page   (starts at 0x800000)
 */ 

   // The memory bus.
   wire [31:0] mem_address; // 24 bits are used internally. The two LSBs are ignored (using word addresses)
   wire  [3:0] mem_wmask;   // mem write mask and strobe /write Legal values are 000,0001,0010,0100,1000,0011,1100,1111
   wire [31:0] mem_rdata;   // processor <- (mem and peripherals) 
   wire [31:0] mem_wdata;   // processor -> (mem and peripherals)
   wire        mem_rstrb;   // mem read strobe. Goes high to initiate memory write.
   wire        mem_rbusy;   // processor <- (mem and peripherals). Stays high until a read transfer is finished.
   wire        mem_wbusy;   // processor <- (mem and peripherals). Stays high until a write transfer is finished.

   wire        mem_wstrb = |mem_wmask; // mem write strobe, goes high to initiate memory write (deduced from wmask)

   // IO bus.
   wire mem_address_is_io  =  mem_address[22];
   wire mem_address_is_ram = !mem_address[22];
      
   reg  [31:0] io_rdata; 
   wire [31:0] io_wdata = mem_wdata;
   wire        io_rstrb = mem_rstrb && mem_address_is_io;
   wire        io_wstrb = mem_wstrb && mem_address_is_io;
   wire [19:0] io_word_address = mem_address[21:2]; // word offset in io page
   wire        io_rbusy; 
   wire        io_wbusy;

   assign      mem_rbusy = io_rbusy;
   assign      mem_wbusy = io_wbusy; 

   wire [19:0] ram_word_address = mem_address[21:2];

// Synthethizing BRAM

   (* no_rw_check *)
   reg [31:0] RAM[0:(`NRV_RAM_SIZE/4)-1];
   reg [31:0] ram_rdata;

   // Initialize the RAM with the generated firmware hex file.
   // The hex file is generated by the bundled elf-2-verilog converter (see TOOLS/FIRMWARE_WORDS_SRC)
   initial begin
      $readmemh("D:/Projects/learn-fpga/blinker_loop.hex",RAM); 
   end

   // The power of YOSYS: it infers BRAM primitives automatically ! (and recognizes
   // masked writes, amazing ...)
   /* verilator lint_off WIDTH */
   always @(posedge clk) begin
      if(mem_address_is_ram) begin
         if(mem_wmask[0]) RAM[ram_word_address][ 7:0 ] <= mem_wdata[ 7:0 ];
         if(mem_wmask[1]) RAM[ram_word_address][15:8 ] <= mem_wdata[15:8 ];
         if(mem_wmask[2]) RAM[ram_word_address][23:16] <= mem_wdata[23:16];
         if(mem_wmask[3]) RAM[ram_word_address][31:24] <= mem_wdata[31:24];	 
      end
      ram_rdata <= RAM[ram_word_address];
   end
   /* verilator lint_on WIDTH */

   assign mem_rdata = mem_address_is_io ? io_rdata : ram_rdata;

/***************************************************************************************************
 *
 * Memory-mapped IO
 * Mapped IO uses "one-hot" addressing, to make decoder
 * simpler (saves a lot of LUTs), as in J1/swapforth,
 * thanks to Matthias Koch(Mecrisp author) for the idea !
 * The included files contains the symbolic constants that
 * determine which device uses which bit.
 */  

`include "HardwareConfig_bits.v"   

/*
 * Devices are components plugged to the IO memory bus.
 * A few words follow in case you want to write your own devices:
 *
 * Each device has one or several register(s). Each register 
 * can be optionally read or/and written.
 * - Each register is selected by a .sel_xxx signal (where xxx
 *   is the name of the register). With the 1-hot encoding that 
 *   I'm using, .sel_xxx is systematically one of the bits of the 
 *   IO word address (it is also possible to write a real
 *   address decoder, at the expense of eating-up a larger 
 *   number of LUTs).
 * - If the device requires wait cycles for writing and/or reading, 
 *   it can have a .wbusy and/or .rbusy signal(s). All the .wbusy
 *   and .rbusy signals of all the devices are ORed at the end of
 *   this file to form the .io_rbusy and .io_wbusy signals.
 * - If the device has read access, then it has a 32-bits .xxx_rdata
 *   signal, that returns 32'b0 if the device is not selected, or the
 *   read data otherwise. All the .xxx_rdata signals of all the devices
 *   are ORed at the end of this file to form the 32-bits io_rdata signal.
 * - Finally, of course, each device is plugged to some pins of the FPGA,
 *   the corresponding signals are in capital letters. 
 */   


/*********************** Hardware configuration ************/
/*
 * Three memory-mapped constant registers that make it easy for
 * client code to query installed RAM and configured devices
 * (this one does not use any pin, of course).
 * Uses some LUTs, a bit stupid, but more comfortable, so that
 * I do not need to change the software on the SDCard each time 
 * I test a different hardware configuration.
 */
`ifdef NRV_IO_HARDWARE_CONFIG   
   wire [31:0] hwconfig_rdata;
   HardwareConfig hwconfig (
      .clk(clk)
     ,.sel_memory(io_word_address[IO_HW_CONFIG_RAM_bit])
     ,.sel_devices(io_word_address[IO_HW_CONFIG_DEVICES_bit])
     ,.sel_cpuinfo(io_word_address[IO_HW_CONFIG_CPUINFO_bit])
     ,.rdata(hwconfig_rdata)
   );
`endif

/*********************** Four LEDs ************************/
`ifdef NRV_IO_LEDS
   wire [31:0] leds_rdata;
   LEDDriver leds (
      .clk(clk)
     ,.rstrb(io_rstrb)
     ,.wstrb(io_wstrb)
     ,.sel(io_word_address[IO_LEDS_bit])
     ,.wdata(io_wdata)
     ,.rdata(leds_rdata)
     ,.LED({D4,D3,D2,D1})
   );
`endif

/********************** SSD1351/SSD1331 oled display ******/
`ifdef NRV_IO_SSD1351_1331
   wire SSD1351_wbusy;
   SSD1351 oled_display (
      .clk(clk)
     ,.RST(oled_RST)
     ,.wstrb(io_wstrb)
     ,.sel_cntl(io_word_address[IO_SSD1351_CNTL_bit])
     ,.sel_cmd(io_word_address[IO_SSD1351_CMD_bit])
     ,.sel_dat(io_word_address[IO_SSD1351_DAT_bit])
     ,.sel_dat16(io_word_address[IO_SSD1351_DAT16_bit])
     ,.wdata(io_wdata)
     ,.wbusy(SSD1351_wbusy)
     ,.DIN(oled_DIN)
     ,.CLK(oled_CLK)
     ,.CS(oled_CS)
     ,.DC(oled_DC)
   );
`endif   

/********************** UART ****************************************/
`ifdef NRV_IO_UART

   // Internal wires to connect IO buffers to UART
   wire RXD_internal;
   wire TXD_internal;

`ifdef ULX3S
   `ifndef BENCH_OR_LINT
     // On the ULX3S, we need to latch RXD, using the latch
     // embedded in the input buffer. If we do not do that,
     // then we unpredictably get garbage on the UART.
     // The two primitives BB (bidirectional three-state buffer)
     // and IFS1P3BX (latch in IO pin) are interpreted by the
     // synthesis tool as an IO cell.
     wire RXD_btw;
     BB RXD_bb(
       .I(1'b0), 
       .O(RXD_btw), 
       .B(RXD), 
       .T(1'b1)
     );
     IFS1P3BX RXD_pin(
       .SCLK(clk),		    
       .D(RXD_btw),
       .Q(RXD_internal),
       .PD(1'b0)		    
     );
     assign TXD = TXD_internal; // For now, do not latch output (but we may need to)
     `define UART_IO_BUFFER
   `endif
 `endif
 
 // For other boards, we directly connect RXD and TXD to the UART (but we may need
 // to latch).
`ifndef UART_IO_BUFFER
   assign RXD_internal = RXD;
   assign TXD = TXD_internal;
`endif

   wire        uart_brk;
   wire [31:0] uart_rdata;
   UART #(
      .NRV_FREQ(`NRV_FREQ)
     ,.NRV_BAUD_RATE(115200)
   ) uart (
      .clk(clk)
     ,.rstrb(io_rstrb)
     ,.wstrb(io_wstrb)
     ,.sel_dat(io_word_address[IO_UART_DAT_bit])
     ,.sel_cntl(io_word_address[IO_UART_CNTL_bit])
     ,.wdata(io_wdata)
     ,.rdata(uart_rdata)
     ,.RXD(RXD_internal)
     ,.TXD(TXD_internal)
     ,.brk(uart_brk)
   );
`else
   wire uart_brk = 1'b0;
`endif

/********** MAX7219 led matrix driver *******************************/
`ifdef NRV_IO_MAX7219
   wire max7219_wbusy;
   MAX7219 max7219 (
      .clk(clk)
     ,.CS(ledmtx_CS)
     ,.wstrb(io_wstrb)
     ,.sel(io_word_address[IO_MAX7219_DAT_bit])
     ,.wdata(io_wdata)
     ,.wbusy(max7219_wbusy)
     ,.DIN(ledmtx_DIN)
     ,.CLK(ledmtx_CLK)
   );
`endif   
   
/********************* SPI SDCard  *********************************/
/*
 * This one has an output register directly wired to the CLK,MOSI,CS_N
 * and an input register directly wired to MISO. The software driver
 * implements the SPI protocol by bit-banging (see FIRMWARE/LIBFEMTORV32/spi_sd.c).
 * One day I'll replace it with a hardware driver... if I have time !
 * ... a generic SPI driver would be good to have also.
 */
`ifdef NRV_IO_SDCARD
   wire [31:0] sdcard_rdata;
   SDCard sdcard (
      .clk(clk)
     ,.rstrb(io_rstrb)
     ,.wstrb(io_wstrb)
     ,.sel(io_word_address[IO_SDCARD_bit])
     ,.wdata(io_wdata)
     ,.rdata(sdcard_rdata)
     ,.CLK(sd_clk)
     ,.MISO(sd_miso)
     ,.MOSI(sd_mosi)
     ,.CS_N(sd_cs_n)
   );
`endif

/********************* Buttons  *************************************/
/*
 * Directly wired to the buttons.
 */
`ifdef NRV_IO_BUTTONS
   wire [31:0] buttons_rdata;
   Buttons buttons_driver (
      .sel(io_word_address[IO_BUTTONS_bit])
     ,.rdata(buttons_rdata)
     ,.BUTTONS(buttons)
   );
`endif
   
/************** io_rdata, io_rbusy and io_wbusy signals *************/

/*
 * io_rdata is latched. Not mandatory, but probably allow higher freq, to be tested.
 */
always @(posedge clk) begin
   io_rdata <= 0
`ifdef NRV_IO_HARDWARE_CONFIG
            | hwconfig_rdata
`endif
`ifdef NRV_IO_LEDS
            | leds_rdata
`endif
`ifdef NRV_IO_UART
            | uart_rdata
`endif
`ifdef NRV_IO_SDCARD
            | sdcard_rdata
`endif
`ifdef NRV_IO_BUTTONS
            | buttons_rdata
`endif
            ;
end

   // For now, we got no device that has
   // blocking reads (SPI flash blocks on
   // write address and waits for read data).
   assign io_rbusy = 0;

   assign io_wbusy = 0
`ifdef NRV_IO_SSD1351_1331
                   | SSD1351_wbusy
`endif
`ifdef NRV_IO_MAX7219
                   | max7219_wbusy
`endif
`ifdef NRV_IO_SPI_FLASH
                   | spi_flash_wbusy
`endif
;

/****************************************************************/
/* And last but not least, the processor                        */

   reg error=1'b0;

  FemtoRV32 #(
      .ADDR_WIDTH(`NRV_ADDR_WIDTH)
     ,.RESET_ADDR(`NRV_RESET_ADDR)
  ) processor (
      .clk(clk)
     ,.mem_addr(mem_address)
     ,.mem_wdata(mem_wdata)
     ,.mem_wmask(mem_wmask)
     ,.mem_rdata(mem_rdata)
     ,.mem_rstrb(mem_rstrb)
     ,.mem_rbusy(mem_rbusy)
     ,.mem_wbusy(mem_wbusy)
`ifdef NRV_INTERRUPTS
     ,.interrupt_request(1'b0)
`endif
     ,.reset(reset && !uart_brk)
   );

`ifdef NRV_IO_LEDS  
   assign D5 = error;
`endif

endmodule


module HardwareConfig (
   input wire 	       clk
  ,input wire 	       sel_memory   // available RAM
  ,input wire 	       sel_devices  // configured devices 
  ,input wire         sel_cpuinfo  // CPU information 	      
  ,output wire [31:0] rdata        // read data
);

`include "HardwareConfig_bits.v"

`ifdef NRV_COUNTER_WIDTH
   localparam counter_width = `NRV_COUNTER_WIDTH;
`else
   localparam counter_width = 32;
`endif   

   
// configured devices
localparam NRV_DEVICES = 0
`ifdef NRV_IO_LEDS
   | (1 << IO_LEDS_bit)
`endif
`ifdef NRV_IO_UART
   | (1 << IO_UART_DAT_bit) | (1 << IO_UART_CNTL_bit)
`endif
`ifdef NRV_IO_SSD1351_1331
   | (1 << IO_SSD1351_CNTL_bit) | (1 << IO_SSD1351_CMD_bit) | (1 << IO_SSD1351_DAT_bit)  
`endif
`ifdef NRV_IO_MAX7219     
   | (1 << IO_MAX7219_DAT_bit) 
`endif
`ifdef NRV_IO_SPI_FLASH
   | (1 << IO_SPI_FLASH_bit)
`endif
`ifdef NRV_MAPPED_SPI_FLASH
   | (1 << IO_MAPPED_SPI_FLASH_bit)
`endif
`ifdef NRV_IO_SDCARD
   | (1 << IO_SDCARD_bit)
`endif
`ifdef NRV_IO_BUTTONS
   | (1 << IO_BUTTONS_bit)
`endif 
`ifdef NRV_IO_FGA
   | (1 << IO_FGA_CNTL_bit) | (1 << IO_FGA_DAT_bit)
`endif
;

   assign rdata = sel_memory  ? `NRV_RAM_SIZE :
                  sel_devices ?  NRV_DEVICES :
                  sel_cpuinfo ? (`NRV_FREQ << 16) | counter_width : 32'b0;

endmodule
